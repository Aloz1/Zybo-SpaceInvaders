----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 24.04.2018 14:18:15
-- Design Name: 
-- Module Name: PSX_Decode_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PSX_Decode_tb is
--  Port ( );
end PSX_Decode_tb;

architecture Behavioral of PSX_Decode_tb is
    constant CLOCK_TICKS  : integer := 400; -- 400 ticks for 250kHz, 14200 ticks for 7kHz
    constant CLOCK_PERIOD : time := 10 ns;
	 
    signal in_clock      : std_logic;
	signal in_reset      : std_logic;
	 
	 
	signal out_done_strb : std_logic;
	signal out_busy      : std_logic;
	signal out_wait_ack  : std_logic;
	signal out_err       : std_logic;
	signal out_data      : std_logic_vector(7 downto 0);
	signal in_atn        : std_logic_vector(1 downto 0);
	signal in_start      : std_logic;
	signal in_cmd        : std_logic_vector(7 downto 0);
	 
	signal out_pin_clock : std_logic;
	signal out_pin_atn   : std_logic_vector(1 downto 0);
	signal in_pin_ack    : std_logic;
	 
	signal out_pin_cmd   : std_logic;
	signal in_pin_data   : std_logic;
begin

     -- Instantiate controller decoder for testing
     PSX_Decode_inst : entity work.PSX_Decode
     generic map (
         C_CLOCK_PERIOD_TICKS => CLOCK_TICKS
     )
     port map (
         s_axi_clock => in_clock,
         s_axi_reset => in_reset,
         
         -- PS control signals
         s_ctrl_done_strb => out_done_strb,
         s_ctrl_busy      => out_busy,
         s_ctrl_wait_ack  => out_wait_ack,
         s_ctrl_err       => out_err,
         s_ctrl_data      => out_data,
         s_ctrl_atn       => in_atn,
         s_ctrl_start     => in_start,
         s_ctrl_cmd       => in_cmd,
         
         -- Control signals
         s_pin_clock => out_pin_clock,
         s_pin_atn   => out_pin_atn,
         s_ack   => in_pin_ack,
         
         -- Command/Data signals
         s_pin_cmd   => out_pin_cmd,
         s_data  => in_pin_data
     );
	 
     -- Heartbeat process
	 process
	 begin
	   in_clock <= '1';
		wait for CLOCK_PERIOD / 2;
		in_clock <= '0';
		wait for CLOCK_PERIOD / 2;
	 end process;
	 
     -- Testcase process
	 process
	 begin
        -- Start by resetting everything
		in_reset    <= '0';
		in_pin_data <= '1';
		in_pin_ack  <= '1';
		in_atn      <= "00";
		in_cmd      <= (others => '0');
		in_start    <= '0';
		
		wait for CLOCK_PERIOD * 5;
		
		in_reset <= '1';
		
		wait for CLOCK_PERIOD * 5;
		
        -- After a couple clock cycles, change ATN
		in_atn <= "10";
		
		wait for CLOCK_PERIOD * 5;
		
        -- Now set CMD (in_start is generated by the AXI interface)
		in_cmd <= x"01";
		in_start   <= '1';
		
        -- Because it's a strobe, it needs to be set back to 0
		wait for CLOCK_PERIOD;
		in_start <= '0';

        -- Bit 0 from PSX
        wait for CLOCK_PERIOD * CLOCK_TICKS - 1;
		in_pin_data <= '0';
		
        -- Bit 1 from PSX
		wait for CLOCK_PERIOD * CLOCK_TICKS * 2;
		in_pin_data <= '1';
		
        -- Bit 2 from PSX
		wait for CLOCK_PERIOD * CLOCK_TICKS * 2;
		in_pin_data <= '0';
		
        -- Bit 3 from PSX
		wait for CLOCK_PERIOD * CLOCK_TICKS * 2;
		in_pin_data <= '1';
		
        -- Bit 4 from PSX
		wait for CLOCK_PERIOD * CLOCK_TICKS * 2;
		in_pin_data <= '0';
		
        -- Bit 5 from PSX
		wait for CLOCK_PERIOD * CLOCK_TICKS * 2;
		in_pin_data <= '1';
		
        -- Bit 6 from PSX
		wait for CLOCK_PERIOD * CLOCK_TICKS * 2;
		in_pin_data <= '0';
		
        -- Bit 7 from PSX
		wait for CLOCK_PERIOD * CLOCK_TICKS * 2;
		in_pin_data <= '1';
		
        -- Send ACK low
		wait for CLOCK_PERIOD * CLOCK_TICKS * 2;
		in_pin_ack  <= '0';
		
        -- Return ACK to high
        wait for CLOCK_PERIOD * CLOCK_TICKS;
		in_pin_ack  <= '1';
		
        -- Reset atn to idle state
		wait for CLOCK_PERIOD * CLOCK_TICKS;
		in_atn <= "11";
		
		wait;
	 end process;
    
end Behavioral;
